-- megafunction wizard: %LPM_DECODE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_DECODE 

-- ============================================================
-- File Name: decode.vhd
-- Megafunction Name(s):
-- 			LPM_DECODE
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.all;

ENTITY decode IS
	PORT
	(
		data		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		eq0		: OUT STD_LOGIC ;
		eq1		: OUT STD_LOGIC ;
		eq10		: OUT STD_LOGIC ;
		eq11		: OUT STD_LOGIC ;
		eq12		: OUT STD_LOGIC ;
		eq13		: OUT STD_LOGIC ;
		eq14		: OUT STD_LOGIC ;
		eq15		: OUT STD_LOGIC ;
		eq16		: OUT STD_LOGIC ;
		eq17		: OUT STD_LOGIC ;
		eq18		: OUT STD_LOGIC ;
		eq19		: OUT STD_LOGIC ;
		eq2		: OUT STD_LOGIC ;
		eq20		: OUT STD_LOGIC ;
		eq21		: OUT STD_LOGIC ;
		eq22		: OUT STD_LOGIC ;
		eq23		: OUT STD_LOGIC ;
		eq24		: OUT STD_LOGIC ;
		eq25		: OUT STD_LOGIC ;
		eq26		: OUT STD_LOGIC ;
		eq27		: OUT STD_LOGIC ;
		eq28		: OUT STD_LOGIC ;
		eq29		: OUT STD_LOGIC ;
		eq3		: OUT STD_LOGIC ;
		eq30		: OUT STD_LOGIC ;
		eq31		: OUT STD_LOGIC ;
		eq32		: OUT STD_LOGIC ;
		eq33		: OUT STD_LOGIC ;
		eq34		: OUT STD_LOGIC ;
		eq35		: OUT STD_LOGIC ;
		eq36		: OUT STD_LOGIC ;
		eq37		: OUT STD_LOGIC ;
		eq38		: OUT STD_LOGIC ;
		eq39		: OUT STD_LOGIC ;
		eq4		: OUT STD_LOGIC ;
		eq40		: OUT STD_LOGIC ;
		eq41		: OUT STD_LOGIC ;
		eq42		: OUT STD_LOGIC ;
		eq43		: OUT STD_LOGIC ;
		eq44		: OUT STD_LOGIC ;
		eq45		: OUT STD_LOGIC ;
		eq46		: OUT STD_LOGIC ;
		eq47		: OUT STD_LOGIC ;
		eq48		: OUT STD_LOGIC ;
		eq49		: OUT STD_LOGIC ;
		eq5		: OUT STD_LOGIC ;
		eq50		: OUT STD_LOGIC ;
		eq51		: OUT STD_LOGIC ;
		eq52		: OUT STD_LOGIC ;
		eq53		: OUT STD_LOGIC ;
		eq54		: OUT STD_LOGIC ;
		eq55		: OUT STD_LOGIC ;
		eq56		: OUT STD_LOGIC ;
		eq57		: OUT STD_LOGIC ;
		eq58		: OUT STD_LOGIC ;
		eq59		: OUT STD_LOGIC ;
		eq6		: OUT STD_LOGIC ;
		eq60		: OUT STD_LOGIC ;
		eq61		: OUT STD_LOGIC ;
		eq62		: OUT STD_LOGIC ;
		eq63		: OUT STD_LOGIC ;
		eq64		: OUT STD_LOGIC ;
		eq65		: OUT STD_LOGIC ;
		eq66		: OUT STD_LOGIC ;
		eq67		: OUT STD_LOGIC ;
		eq68		: OUT STD_LOGIC ;
		eq69		: OUT STD_LOGIC ;
		eq7		: OUT STD_LOGIC ;
		eq70		: OUT STD_LOGIC ;
		eq8		: OUT STD_LOGIC ;
		eq9		: OUT STD_LOGIC 
	);
END decode;


ARCHITECTURE SYN OF decode IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC ;
	SIGNAL sub_wire3	: STD_LOGIC ;
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC ;
	SIGNAL sub_wire6	: STD_LOGIC ;
	SIGNAL sub_wire7	: STD_LOGIC ;
	SIGNAL sub_wire8	: STD_LOGIC ;
	SIGNAL sub_wire9	: STD_LOGIC ;
	SIGNAL sub_wire10	: STD_LOGIC ;
	SIGNAL sub_wire11	: STD_LOGIC ;
	SIGNAL sub_wire12	: STD_LOGIC ;
	SIGNAL sub_wire13	: STD_LOGIC ;
	SIGNAL sub_wire14	: STD_LOGIC ;
	SIGNAL sub_wire15	: STD_LOGIC ;
	SIGNAL sub_wire16	: STD_LOGIC ;
	SIGNAL sub_wire17	: STD_LOGIC ;
	SIGNAL sub_wire18	: STD_LOGIC ;
	SIGNAL sub_wire19	: STD_LOGIC ;
	SIGNAL sub_wire20	: STD_LOGIC ;
	SIGNAL sub_wire21	: STD_LOGIC ;
	SIGNAL sub_wire22	: STD_LOGIC ;
	SIGNAL sub_wire23	: STD_LOGIC ;
	SIGNAL sub_wire24	: STD_LOGIC ;
	SIGNAL sub_wire25	: STD_LOGIC ;
	SIGNAL sub_wire26	: STD_LOGIC ;
	SIGNAL sub_wire27	: STD_LOGIC ;
	SIGNAL sub_wire28	: STD_LOGIC ;
	SIGNAL sub_wire29	: STD_LOGIC ;
	SIGNAL sub_wire30	: STD_LOGIC ;
	SIGNAL sub_wire31	: STD_LOGIC ;
	SIGNAL sub_wire32	: STD_LOGIC ;
	SIGNAL sub_wire33	: STD_LOGIC ;
	SIGNAL sub_wire34	: STD_LOGIC ;
	SIGNAL sub_wire35	: STD_LOGIC ;
	SIGNAL sub_wire36	: STD_LOGIC ;
	SIGNAL sub_wire37	: STD_LOGIC ;
	SIGNAL sub_wire38	: STD_LOGIC ;
	SIGNAL sub_wire39	: STD_LOGIC ;
	SIGNAL sub_wire40	: STD_LOGIC ;
	SIGNAL sub_wire41	: STD_LOGIC ;
	SIGNAL sub_wire42	: STD_LOGIC ;
	SIGNAL sub_wire43	: STD_LOGIC ;
	SIGNAL sub_wire44	: STD_LOGIC ;
	SIGNAL sub_wire45	: STD_LOGIC ;
	SIGNAL sub_wire46	: STD_LOGIC ;
	SIGNAL sub_wire47	: STD_LOGIC ;
	SIGNAL sub_wire48	: STD_LOGIC ;
	SIGNAL sub_wire49	: STD_LOGIC ;
	SIGNAL sub_wire50	: STD_LOGIC ;
	SIGNAL sub_wire51	: STD_LOGIC ;
	SIGNAL sub_wire52	: STD_LOGIC ;
	SIGNAL sub_wire53	: STD_LOGIC ;
	SIGNAL sub_wire54	: STD_LOGIC ;
	SIGNAL sub_wire55	: STD_LOGIC ;
	SIGNAL sub_wire56	: STD_LOGIC ;
	SIGNAL sub_wire57	: STD_LOGIC ;
	SIGNAL sub_wire58	: STD_LOGIC ;
	SIGNAL sub_wire59	: STD_LOGIC ;
	SIGNAL sub_wire60	: STD_LOGIC ;
	SIGNAL sub_wire61	: STD_LOGIC ;
	SIGNAL sub_wire62	: STD_LOGIC ;
	SIGNAL sub_wire63	: STD_LOGIC ;
	SIGNAL sub_wire64	: STD_LOGIC ;
	SIGNAL sub_wire65	: STD_LOGIC ;
	SIGNAL sub_wire66	: STD_LOGIC ;
	SIGNAL sub_wire67	: STD_LOGIC ;
	SIGNAL sub_wire68	: STD_LOGIC ;
	SIGNAL sub_wire69	: STD_LOGIC ;
	SIGNAL sub_wire70	: STD_LOGIC ;
	SIGNAL sub_wire71	: STD_LOGIC ;



	COMPONENT lpm_decode
	GENERIC (
		lpm_decodes		: NATURAL;
		lpm_type		: STRING;
		lpm_width		: NATURAL
	);
	PORT (
			data	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			eq	: OUT STD_LOGIC_VECTOR (255 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	sub_wire71    <= sub_wire0(65);
	sub_wire70    <= sub_wire0(47);
	sub_wire69    <= sub_wire0(29);
	sub_wire68    <= sub_wire0(64);
	sub_wire67    <= sub_wire0(46);
	sub_wire66    <= sub_wire0(28);
	sub_wire65    <= sub_wire0(9);
	sub_wire64    <= sub_wire0(63);
	sub_wire63    <= sub_wire0(54);
	sub_wire62    <= sub_wire0(45);
	sub_wire61    <= sub_wire0(36);
	sub_wire60    <= sub_wire0(27);
	sub_wire59    <= sub_wire0(18);
	sub_wire58    <= sub_wire0(8);
	sub_wire57    <= sub_wire0(62);
	sub_wire56    <= sub_wire0(53);
	sub_wire55    <= sub_wire0(44);
	sub_wire54    <= sub_wire0(35);
	sub_wire53    <= sub_wire0(26);
	sub_wire52    <= sub_wire0(17);
	sub_wire51    <= sub_wire0(70);
	sub_wire50    <= sub_wire0(7);
	sub_wire49    <= sub_wire0(61);
	sub_wire48    <= sub_wire0(52);
	sub_wire47    <= sub_wire0(43);
	sub_wire46    <= sub_wire0(34);
	sub_wire45    <= sub_wire0(25);
	sub_wire44    <= sub_wire0(16);
	sub_wire43    <= sub_wire0(60);
	sub_wire42    <= sub_wire0(6);
	sub_wire41    <= sub_wire0(51);
	sub_wire40    <= sub_wire0(42);
	sub_wire39    <= sub_wire0(33);
	sub_wire38    <= sub_wire0(24);
	sub_wire37    <= sub_wire0(15);
	sub_wire36    <= sub_wire0(50);
	sub_wire35    <= sub_wire0(5);
	sub_wire34    <= sub_wire0(41);
	sub_wire33    <= sub_wire0(32);
	sub_wire32    <= sub_wire0(23);
	sub_wire31    <= sub_wire0(14);
	sub_wire30    <= sub_wire0(40);
	sub_wire29    <= sub_wire0(4);
	sub_wire28    <= sub_wire0(31);
	sub_wire27    <= sub_wire0(22);
	sub_wire26    <= sub_wire0(13);
	sub_wire25    <= sub_wire0(30);
	sub_wire24    <= sub_wire0(3);
	sub_wire23    <= sub_wire0(21);
	sub_wire22    <= sub_wire0(12);
	sub_wire21    <= sub_wire0(20);
	sub_wire20    <= sub_wire0(2);
	sub_wire19    <= sub_wire0(11);
	sub_wire18    <= sub_wire0(10);
	sub_wire17    <= sub_wire0(1);
	sub_wire16    <= sub_wire0(0);
	sub_wire15    <= sub_wire0(69);
	sub_wire14    <= sub_wire0(68);
	sub_wire13    <= sub_wire0(59);
	sub_wire12    <= sub_wire0(67);
	sub_wire11    <= sub_wire0(58);
	sub_wire10    <= sub_wire0(49);
	sub_wire9    <= sub_wire0(66);
	sub_wire8    <= sub_wire0(57);
	sub_wire7    <= sub_wire0(48);
	sub_wire6    <= sub_wire0(39);
	sub_wire5    <= sub_wire0(56);
	sub_wire4    <= sub_wire0(38);
	sub_wire3    <= sub_wire0(55);
	sub_wire2    <= sub_wire0(37);
	sub_wire1    <= sub_wire0(19);
	eq19    <= sub_wire1;
	eq37    <= sub_wire2;
	eq55    <= sub_wire3;
	eq38    <= sub_wire4;
	eq56    <= sub_wire5;
	eq39    <= sub_wire6;
	eq48    <= sub_wire7;
	eq57    <= sub_wire8;
	eq66    <= sub_wire9;
	eq49    <= sub_wire10;
	eq58    <= sub_wire11;
	eq67    <= sub_wire12;
	eq59    <= sub_wire13;
	eq68    <= sub_wire14;
	eq69    <= sub_wire15;
	eq0    <= sub_wire16;
	eq1    <= sub_wire17;
	eq10    <= sub_wire18;
	eq11    <= sub_wire19;
	eq2    <= sub_wire20;
	eq20    <= sub_wire21;
	eq12    <= sub_wire22;
	eq21    <= sub_wire23;
	eq3    <= sub_wire24;
	eq30    <= sub_wire25;
	eq13    <= sub_wire26;
	eq22    <= sub_wire27;
	eq31    <= sub_wire28;
	eq4    <= sub_wire29;
	eq40    <= sub_wire30;
	eq14    <= sub_wire31;
	eq23    <= sub_wire32;
	eq32    <= sub_wire33;
	eq41    <= sub_wire34;
	eq5    <= sub_wire35;
	eq50    <= sub_wire36;
	eq15    <= sub_wire37;
	eq24    <= sub_wire38;
	eq33    <= sub_wire39;
	eq42    <= sub_wire40;
	eq51    <= sub_wire41;
	eq6    <= sub_wire42;
	eq60    <= sub_wire43;
	eq16    <= sub_wire44;
	eq25    <= sub_wire45;
	eq34    <= sub_wire46;
	eq43    <= sub_wire47;
	eq52    <= sub_wire48;
	eq61    <= sub_wire49;
	eq7    <= sub_wire50;
	eq70    <= sub_wire51;
	eq17    <= sub_wire52;
	eq26    <= sub_wire53;
	eq35    <= sub_wire54;
	eq44    <= sub_wire55;
	eq53    <= sub_wire56;
	eq62    <= sub_wire57;
	eq8    <= sub_wire58;
	eq18    <= sub_wire59;
	eq27    <= sub_wire60;
	eq36    <= sub_wire61;
	eq45    <= sub_wire62;
	eq54    <= sub_wire63;
	eq63    <= sub_wire64;
	eq9    <= sub_wire65;
	eq28    <= sub_wire66;
	eq46    <= sub_wire67;
	eq64    <= sub_wire68;
	eq29    <= sub_wire69;
	eq47    <= sub_wire70;
	eq65    <= sub_wire71;

	LPM_DECODE_component : LPM_DECODE
	GENERIC MAP (
		lpm_decodes => 256,
		lpm_type => "LPM_DECODE",
		lpm_width => 8
	)
	PORT MAP (
		data => data,
		eq => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: BaseDec NUMERIC "1"
-- Retrieval info: PRIVATE: EnableInput NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
-- Retrieval info: PRIVATE: Latency NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: aclr NUMERIC "0"
-- Retrieval info: PRIVATE: clken NUMERIC "0"
-- Retrieval info: PRIVATE: eq0 NUMERIC "1"
-- Retrieval info: PRIVATE: eq1 NUMERIC "1"
-- Retrieval info: PRIVATE: eq10 NUMERIC "1"
-- Retrieval info: PRIVATE: eq100 NUMERIC "0"
-- Retrieval info: PRIVATE: eq101 NUMERIC "0"
-- Retrieval info: PRIVATE: eq102 NUMERIC "0"
-- Retrieval info: PRIVATE: eq103 NUMERIC "0"
-- Retrieval info: PRIVATE: eq104 NUMERIC "0"
-- Retrieval info: PRIVATE: eq105 NUMERIC "0"
-- Retrieval info: PRIVATE: eq106 NUMERIC "0"
-- Retrieval info: PRIVATE: eq107 NUMERIC "0"
-- Retrieval info: PRIVATE: eq108 NUMERIC "0"
-- Retrieval info: PRIVATE: eq109 NUMERIC "0"
-- Retrieval info: PRIVATE: eq11 NUMERIC "1"
-- Retrieval info: PRIVATE: eq110 NUMERIC "0"
-- Retrieval info: PRIVATE: eq111 NUMERIC "0"
-- Retrieval info: PRIVATE: eq112 NUMERIC "0"
-- Retrieval info: PRIVATE: eq113 NUMERIC "0"
-- Retrieval info: PRIVATE: eq114 NUMERIC "0"
-- Retrieval info: PRIVATE: eq115 NUMERIC "0"
-- Retrieval info: PRIVATE: eq116 NUMERIC "0"
-- Retrieval info: PRIVATE: eq117 NUMERIC "0"
-- Retrieval info: PRIVATE: eq118 NUMERIC "0"
-- Retrieval info: PRIVATE: eq119 NUMERIC "0"
-- Retrieval info: PRIVATE: eq12 NUMERIC "1"
-- Retrieval info: PRIVATE: eq120 NUMERIC "0"
-- Retrieval info: PRIVATE: eq121 NUMERIC "0"
-- Retrieval info: PRIVATE: eq122 NUMERIC "0"
-- Retrieval info: PRIVATE: eq123 NUMERIC "0"
-- Retrieval info: PRIVATE: eq124 NUMERIC "0"
-- Retrieval info: PRIVATE: eq125 NUMERIC "0"
-- Retrieval info: PRIVATE: eq126 NUMERIC "0"
-- Retrieval info: PRIVATE: eq127 NUMERIC "0"
-- Retrieval info: PRIVATE: eq128 NUMERIC "0"
-- Retrieval info: PRIVATE: eq129 NUMERIC "0"
-- Retrieval info: PRIVATE: eq13 NUMERIC "1"
-- Retrieval info: PRIVATE: eq130 NUMERIC "0"
-- Retrieval info: PRIVATE: eq131 NUMERIC "0"
-- Retrieval info: PRIVATE: eq132 NUMERIC "0"
-- Retrieval info: PRIVATE: eq133 NUMERIC "0"
-- Retrieval info: PRIVATE: eq134 NUMERIC "0"
-- Retrieval info: PRIVATE: eq135 NUMERIC "0"
-- Retrieval info: PRIVATE: eq136 NUMERIC "0"
-- Retrieval info: PRIVATE: eq137 NUMERIC "0"
-- Retrieval info: PRIVATE: eq138 NUMERIC "0"
-- Retrieval info: PRIVATE: eq139 NUMERIC "0"
-- Retrieval info: PRIVATE: eq14 NUMERIC "1"
-- Retrieval info: PRIVATE: eq140 NUMERIC "0"
-- Retrieval info: PRIVATE: eq141 NUMERIC "0"
-- Retrieval info: PRIVATE: eq142 NUMERIC "0"
-- Retrieval info: PRIVATE: eq143 NUMERIC "0"
-- Retrieval info: PRIVATE: eq144 NUMERIC "0"
-- Retrieval info: PRIVATE: eq145 NUMERIC "0"
-- Retrieval info: PRIVATE: eq146 NUMERIC "0"
-- Retrieval info: PRIVATE: eq147 NUMERIC "0"
-- Retrieval info: PRIVATE: eq148 NUMERIC "0"
-- Retrieval info: PRIVATE: eq149 NUMERIC "0"
-- Retrieval info: PRIVATE: eq15 NUMERIC "1"
-- Retrieval info: PRIVATE: eq150 NUMERIC "0"
-- Retrieval info: PRIVATE: eq151 NUMERIC "0"
-- Retrieval info: PRIVATE: eq152 NUMERIC "0"
-- Retrieval info: PRIVATE: eq153 NUMERIC "0"
-- Retrieval info: PRIVATE: eq154 NUMERIC "0"
-- Retrieval info: PRIVATE: eq155 NUMERIC "0"
-- Retrieval info: PRIVATE: eq156 NUMERIC "0"
-- Retrieval info: PRIVATE: eq157 NUMERIC "0"
-- Retrieval info: PRIVATE: eq158 NUMERIC "0"
-- Retrieval info: PRIVATE: eq159 NUMERIC "0"
-- Retrieval info: PRIVATE: eq16 NUMERIC "1"
-- Retrieval info: PRIVATE: eq160 NUMERIC "0"
-- Retrieval info: PRIVATE: eq161 NUMERIC "0"
-- Retrieval info: PRIVATE: eq162 NUMERIC "0"
-- Retrieval info: PRIVATE: eq163 NUMERIC "0"
-- Retrieval info: PRIVATE: eq164 NUMERIC "0"
-- Retrieval info: PRIVATE: eq165 NUMERIC "0"
-- Retrieval info: PRIVATE: eq166 NUMERIC "0"
-- Retrieval info: PRIVATE: eq167 NUMERIC "0"
-- Retrieval info: PRIVATE: eq168 NUMERIC "0"
-- Retrieval info: PRIVATE: eq169 NUMERIC "0"
-- Retrieval info: PRIVATE: eq17 NUMERIC "1"
-- Retrieval info: PRIVATE: eq170 NUMERIC "0"
-- Retrieval info: PRIVATE: eq171 NUMERIC "0"
-- Retrieval info: PRIVATE: eq172 NUMERIC "0"
-- Retrieval info: PRIVATE: eq173 NUMERIC "0"
-- Retrieval info: PRIVATE: eq174 NUMERIC "0"
-- Retrieval info: PRIVATE: eq175 NUMERIC "0"
-- Retrieval info: PRIVATE: eq176 NUMERIC "0"
-- Retrieval info: PRIVATE: eq177 NUMERIC "0"
-- Retrieval info: PRIVATE: eq178 NUMERIC "0"
-- Retrieval info: PRIVATE: eq179 NUMERIC "0"
-- Retrieval info: PRIVATE: eq18 NUMERIC "1"
-- Retrieval info: PRIVATE: eq180 NUMERIC "0"
-- Retrieval info: PRIVATE: eq181 NUMERIC "0"
-- Retrieval info: PRIVATE: eq182 NUMERIC "0"
-- Retrieval info: PRIVATE: eq183 NUMERIC "0"
-- Retrieval info: PRIVATE: eq184 NUMERIC "0"
-- Retrieval info: PRIVATE: eq185 NUMERIC "0"
-- Retrieval info: PRIVATE: eq186 NUMERIC "0"
-- Retrieval info: PRIVATE: eq187 NUMERIC "0"
-- Retrieval info: PRIVATE: eq188 NUMERIC "0"
-- Retrieval info: PRIVATE: eq189 NUMERIC "0"
-- Retrieval info: PRIVATE: eq19 NUMERIC "1"
-- Retrieval info: PRIVATE: eq190 NUMERIC "0"
-- Retrieval info: PRIVATE: eq191 NUMERIC "0"
-- Retrieval info: PRIVATE: eq192 NUMERIC "0"
-- Retrieval info: PRIVATE: eq193 NUMERIC "0"
-- Retrieval info: PRIVATE: eq194 NUMERIC "0"
-- Retrieval info: PRIVATE: eq195 NUMERIC "0"
-- Retrieval info: PRIVATE: eq196 NUMERIC "0"
-- Retrieval info: PRIVATE: eq197 NUMERIC "0"
-- Retrieval info: PRIVATE: eq198 NUMERIC "0"
-- Retrieval info: PRIVATE: eq199 NUMERIC "0"
-- Retrieval info: PRIVATE: eq2 NUMERIC "1"
-- Retrieval info: PRIVATE: eq20 NUMERIC "1"
-- Retrieval info: PRIVATE: eq200 NUMERIC "0"
-- Retrieval info: PRIVATE: eq201 NUMERIC "0"
-- Retrieval info: PRIVATE: eq202 NUMERIC "0"
-- Retrieval info: PRIVATE: eq203 NUMERIC "0"
-- Retrieval info: PRIVATE: eq204 NUMERIC "0"
-- Retrieval info: PRIVATE: eq205 NUMERIC "0"
-- Retrieval info: PRIVATE: eq206 NUMERIC "0"
-- Retrieval info: PRIVATE: eq207 NUMERIC "0"
-- Retrieval info: PRIVATE: eq208 NUMERIC "0"
-- Retrieval info: PRIVATE: eq209 NUMERIC "0"
-- Retrieval info: PRIVATE: eq21 NUMERIC "1"
-- Retrieval info: PRIVATE: eq210 NUMERIC "0"
-- Retrieval info: PRIVATE: eq211 NUMERIC "0"
-- Retrieval info: PRIVATE: eq212 NUMERIC "0"
-- Retrieval info: PRIVATE: eq213 NUMERIC "0"
-- Retrieval info: PRIVATE: eq214 NUMERIC "0"
-- Retrieval info: PRIVATE: eq215 NUMERIC "0"
-- Retrieval info: PRIVATE: eq216 NUMERIC "0"
-- Retrieval info: PRIVATE: eq217 NUMERIC "0"
-- Retrieval info: PRIVATE: eq218 NUMERIC "0"
-- Retrieval info: PRIVATE: eq219 NUMERIC "0"
-- Retrieval info: PRIVATE: eq22 NUMERIC "1"
-- Retrieval info: PRIVATE: eq220 NUMERIC "0"
-- Retrieval info: PRIVATE: eq221 NUMERIC "0"
-- Retrieval info: PRIVATE: eq222 NUMERIC "0"
-- Retrieval info: PRIVATE: eq223 NUMERIC "0"
-- Retrieval info: PRIVATE: eq224 NUMERIC "0"
-- Retrieval info: PRIVATE: eq225 NUMERIC "0"
-- Retrieval info: PRIVATE: eq226 NUMERIC "0"
-- Retrieval info: PRIVATE: eq227 NUMERIC "0"
-- Retrieval info: PRIVATE: eq228 NUMERIC "0"
-- Retrieval info: PRIVATE: eq229 NUMERIC "0"
-- Retrieval info: PRIVATE: eq23 NUMERIC "1"
-- Retrieval info: PRIVATE: eq230 NUMERIC "0"
-- Retrieval info: PRIVATE: eq231 NUMERIC "0"
-- Retrieval info: PRIVATE: eq232 NUMERIC "0"
-- Retrieval info: PRIVATE: eq233 NUMERIC "0"
-- Retrieval info: PRIVATE: eq234 NUMERIC "0"
-- Retrieval info: PRIVATE: eq235 NUMERIC "0"
-- Retrieval info: PRIVATE: eq236 NUMERIC "0"
-- Retrieval info: PRIVATE: eq237 NUMERIC "0"
-- Retrieval info: PRIVATE: eq238 NUMERIC "0"
-- Retrieval info: PRIVATE: eq239 NUMERIC "0"
-- Retrieval info: PRIVATE: eq24 NUMERIC "1"
-- Retrieval info: PRIVATE: eq240 NUMERIC "0"
-- Retrieval info: PRIVATE: eq241 NUMERIC "0"
-- Retrieval info: PRIVATE: eq242 NUMERIC "0"
-- Retrieval info: PRIVATE: eq243 NUMERIC "0"
-- Retrieval info: PRIVATE: eq244 NUMERIC "0"
-- Retrieval info: PRIVATE: eq245 NUMERIC "0"
-- Retrieval info: PRIVATE: eq246 NUMERIC "0"
-- Retrieval info: PRIVATE: eq247 NUMERIC "0"
-- Retrieval info: PRIVATE: eq248 NUMERIC "0"
-- Retrieval info: PRIVATE: eq249 NUMERIC "0"
-- Retrieval info: PRIVATE: eq25 NUMERIC "1"
-- Retrieval info: PRIVATE: eq250 NUMERIC "0"
-- Retrieval info: PRIVATE: eq251 NUMERIC "0"
-- Retrieval info: PRIVATE: eq252 NUMERIC "0"
-- Retrieval info: PRIVATE: eq253 NUMERIC "0"
-- Retrieval info: PRIVATE: eq254 NUMERIC "0"
-- Retrieval info: PRIVATE: eq255 NUMERIC "0"
-- Retrieval info: PRIVATE: eq26 NUMERIC "1"
-- Retrieval info: PRIVATE: eq27 NUMERIC "1"
-- Retrieval info: PRIVATE: eq28 NUMERIC "1"
-- Retrieval info: PRIVATE: eq29 NUMERIC "1"
-- Retrieval info: PRIVATE: eq3 NUMERIC "1"
-- Retrieval info: PRIVATE: eq30 NUMERIC "1"
-- Retrieval info: PRIVATE: eq31 NUMERIC "1"
-- Retrieval info: PRIVATE: eq32 NUMERIC "1"
-- Retrieval info: PRIVATE: eq33 NUMERIC "1"
-- Retrieval info: PRIVATE: eq34 NUMERIC "1"
-- Retrieval info: PRIVATE: eq35 NUMERIC "1"
-- Retrieval info: PRIVATE: eq36 NUMERIC "1"
-- Retrieval info: PRIVATE: eq37 NUMERIC "1"
-- Retrieval info: PRIVATE: eq38 NUMERIC "1"
-- Retrieval info: PRIVATE: eq39 NUMERIC "1"
-- Retrieval info: PRIVATE: eq4 NUMERIC "1"
-- Retrieval info: PRIVATE: eq40 NUMERIC "1"
-- Retrieval info: PRIVATE: eq41 NUMERIC "1"
-- Retrieval info: PRIVATE: eq42 NUMERIC "1"
-- Retrieval info: PRIVATE: eq43 NUMERIC "1"
-- Retrieval info: PRIVATE: eq44 NUMERIC "1"
-- Retrieval info: PRIVATE: eq45 NUMERIC "1"
-- Retrieval info: PRIVATE: eq46 NUMERIC "1"
-- Retrieval info: PRIVATE: eq47 NUMERIC "1"
-- Retrieval info: PRIVATE: eq48 NUMERIC "1"
-- Retrieval info: PRIVATE: eq49 NUMERIC "1"
-- Retrieval info: PRIVATE: eq5 NUMERIC "1"
-- Retrieval info: PRIVATE: eq50 NUMERIC "1"
-- Retrieval info: PRIVATE: eq51 NUMERIC "1"
-- Retrieval info: PRIVATE: eq52 NUMERIC "1"
-- Retrieval info: PRIVATE: eq53 NUMERIC "1"
-- Retrieval info: PRIVATE: eq54 NUMERIC "1"
-- Retrieval info: PRIVATE: eq55 NUMERIC "1"
-- Retrieval info: PRIVATE: eq56 NUMERIC "1"
-- Retrieval info: PRIVATE: eq57 NUMERIC "1"
-- Retrieval info: PRIVATE: eq58 NUMERIC "1"
-- Retrieval info: PRIVATE: eq59 NUMERIC "1"
-- Retrieval info: PRIVATE: eq6 NUMERIC "1"
-- Retrieval info: PRIVATE: eq60 NUMERIC "1"
-- Retrieval info: PRIVATE: eq61 NUMERIC "1"
-- Retrieval info: PRIVATE: eq62 NUMERIC "1"
-- Retrieval info: PRIVATE: eq63 NUMERIC "1"
-- Retrieval info: PRIVATE: eq64 NUMERIC "1"
-- Retrieval info: PRIVATE: eq65 NUMERIC "1"
-- Retrieval info: PRIVATE: eq66 NUMERIC "1"
-- Retrieval info: PRIVATE: eq67 NUMERIC "1"
-- Retrieval info: PRIVATE: eq68 NUMERIC "1"
-- Retrieval info: PRIVATE: eq69 NUMERIC "1"
-- Retrieval info: PRIVATE: eq7 NUMERIC "1"
-- Retrieval info: PRIVATE: eq70 NUMERIC "1"
-- Retrieval info: PRIVATE: eq71 NUMERIC "0"
-- Retrieval info: PRIVATE: eq72 NUMERIC "0"
-- Retrieval info: PRIVATE: eq73 NUMERIC "0"
-- Retrieval info: PRIVATE: eq74 NUMERIC "0"
-- Retrieval info: PRIVATE: eq75 NUMERIC "0"
-- Retrieval info: PRIVATE: eq76 NUMERIC "0"
-- Retrieval info: PRIVATE: eq77 NUMERIC "0"
-- Retrieval info: PRIVATE: eq78 NUMERIC "0"
-- Retrieval info: PRIVATE: eq79 NUMERIC "0"
-- Retrieval info: PRIVATE: eq8 NUMERIC "1"
-- Retrieval info: PRIVATE: eq80 NUMERIC "0"
-- Retrieval info: PRIVATE: eq81 NUMERIC "0"
-- Retrieval info: PRIVATE: eq82 NUMERIC "0"
-- Retrieval info: PRIVATE: eq83 NUMERIC "0"
-- Retrieval info: PRIVATE: eq84 NUMERIC "0"
-- Retrieval info: PRIVATE: eq85 NUMERIC "0"
-- Retrieval info: PRIVATE: eq86 NUMERIC "0"
-- Retrieval info: PRIVATE: eq87 NUMERIC "0"
-- Retrieval info: PRIVATE: eq88 NUMERIC "0"
-- Retrieval info: PRIVATE: eq89 NUMERIC "0"
-- Retrieval info: PRIVATE: eq9 NUMERIC "1"
-- Retrieval info: PRIVATE: eq90 NUMERIC "0"
-- Retrieval info: PRIVATE: eq91 NUMERIC "0"
-- Retrieval info: PRIVATE: eq92 NUMERIC "0"
-- Retrieval info: PRIVATE: eq93 NUMERIC "0"
-- Retrieval info: PRIVATE: eq94 NUMERIC "0"
-- Retrieval info: PRIVATE: eq95 NUMERIC "0"
-- Retrieval info: PRIVATE: eq96 NUMERIC "0"
-- Retrieval info: PRIVATE: eq97 NUMERIC "0"
-- Retrieval info: PRIVATE: eq98 NUMERIC "0"
-- Retrieval info: PRIVATE: eq99 NUMERIC "0"
-- Retrieval info: PRIVATE: nBit NUMERIC "8"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_DECODES NUMERIC "256"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DECODE"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "8"
-- Retrieval info: USED_PORT: @eq 0 0 256 0 OUTPUT NODEFVAL "@eq[255..0]"
-- Retrieval info: USED_PORT: data 0 0 8 0 INPUT NODEFVAL "data[7..0]"
-- Retrieval info: USED_PORT: eq0 0 0 0 0 OUTPUT NODEFVAL "eq0"
-- Retrieval info: USED_PORT: eq1 0 0 0 0 OUTPUT NODEFVAL "eq1"
-- Retrieval info: USED_PORT: eq10 0 0 0 0 OUTPUT NODEFVAL "eq10"
-- Retrieval info: USED_PORT: eq11 0 0 0 0 OUTPUT NODEFVAL "eq11"
-- Retrieval info: USED_PORT: eq12 0 0 0 0 OUTPUT NODEFVAL "eq12"
-- Retrieval info: USED_PORT: eq13 0 0 0 0 OUTPUT NODEFVAL "eq13"
-- Retrieval info: USED_PORT: eq14 0 0 0 0 OUTPUT NODEFVAL "eq14"
-- Retrieval info: USED_PORT: eq15 0 0 0 0 OUTPUT NODEFVAL "eq15"
-- Retrieval info: USED_PORT: eq16 0 0 0 0 OUTPUT NODEFVAL "eq16"
-- Retrieval info: USED_PORT: eq17 0 0 0 0 OUTPUT NODEFVAL "eq17"
-- Retrieval info: USED_PORT: eq18 0 0 0 0 OUTPUT NODEFVAL "eq18"
-- Retrieval info: USED_PORT: eq19 0 0 0 0 OUTPUT NODEFVAL "eq19"
-- Retrieval info: USED_PORT: eq2 0 0 0 0 OUTPUT NODEFVAL "eq2"
-- Retrieval info: USED_PORT: eq20 0 0 0 0 OUTPUT NODEFVAL "eq20"
-- Retrieval info: USED_PORT: eq21 0 0 0 0 OUTPUT NODEFVAL "eq21"
-- Retrieval info: USED_PORT: eq22 0 0 0 0 OUTPUT NODEFVAL "eq22"
-- Retrieval info: USED_PORT: eq23 0 0 0 0 OUTPUT NODEFVAL "eq23"
-- Retrieval info: USED_PORT: eq24 0 0 0 0 OUTPUT NODEFVAL "eq24"
-- Retrieval info: USED_PORT: eq25 0 0 0 0 OUTPUT NODEFVAL "eq25"
-- Retrieval info: USED_PORT: eq26 0 0 0 0 OUTPUT NODEFVAL "eq26"
-- Retrieval info: USED_PORT: eq27 0 0 0 0 OUTPUT NODEFVAL "eq27"
-- Retrieval info: USED_PORT: eq28 0 0 0 0 OUTPUT NODEFVAL "eq28"
-- Retrieval info: USED_PORT: eq29 0 0 0 0 OUTPUT NODEFVAL "eq29"
-- Retrieval info: USED_PORT: eq3 0 0 0 0 OUTPUT NODEFVAL "eq3"
-- Retrieval info: USED_PORT: eq30 0 0 0 0 OUTPUT NODEFVAL "eq30"
-- Retrieval info: USED_PORT: eq31 0 0 0 0 OUTPUT NODEFVAL "eq31"
-- Retrieval info: USED_PORT: eq32 0 0 0 0 OUTPUT NODEFVAL "eq32"
-- Retrieval info: USED_PORT: eq33 0 0 0 0 OUTPUT NODEFVAL "eq33"
-- Retrieval info: USED_PORT: eq34 0 0 0 0 OUTPUT NODEFVAL "eq34"
-- Retrieval info: USED_PORT: eq35 0 0 0 0 OUTPUT NODEFVAL "eq35"
-- Retrieval info: USED_PORT: eq36 0 0 0 0 OUTPUT NODEFVAL "eq36"
-- Retrieval info: USED_PORT: eq37 0 0 0 0 OUTPUT NODEFVAL "eq37"
-- Retrieval info: USED_PORT: eq38 0 0 0 0 OUTPUT NODEFVAL "eq38"
-- Retrieval info: USED_PORT: eq39 0 0 0 0 OUTPUT NODEFVAL "eq39"
-- Retrieval info: USED_PORT: eq4 0 0 0 0 OUTPUT NODEFVAL "eq4"
-- Retrieval info: USED_PORT: eq40 0 0 0 0 OUTPUT NODEFVAL "eq40"
-- Retrieval info: USED_PORT: eq41 0 0 0 0 OUTPUT NODEFVAL "eq41"
-- Retrieval info: USED_PORT: eq42 0 0 0 0 OUTPUT NODEFVAL "eq42"
-- Retrieval info: USED_PORT: eq43 0 0 0 0 OUTPUT NODEFVAL "eq43"
-- Retrieval info: USED_PORT: eq44 0 0 0 0 OUTPUT NODEFVAL "eq44"
-- Retrieval info: USED_PORT: eq45 0 0 0 0 OUTPUT NODEFVAL "eq45"
-- Retrieval info: USED_PORT: eq46 0 0 0 0 OUTPUT NODEFVAL "eq46"
-- Retrieval info: USED_PORT: eq47 0 0 0 0 OUTPUT NODEFVAL "eq47"
-- Retrieval info: USED_PORT: eq48 0 0 0 0 OUTPUT NODEFVAL "eq48"
-- Retrieval info: USED_PORT: eq49 0 0 0 0 OUTPUT NODEFVAL "eq49"
-- Retrieval info: USED_PORT: eq5 0 0 0 0 OUTPUT NODEFVAL "eq5"
-- Retrieval info: USED_PORT: eq50 0 0 0 0 OUTPUT NODEFVAL "eq50"
-- Retrieval info: USED_PORT: eq51 0 0 0 0 OUTPUT NODEFVAL "eq51"
-- Retrieval info: USED_PORT: eq52 0 0 0 0 OUTPUT NODEFVAL "eq52"
-- Retrieval info: USED_PORT: eq53 0 0 0 0 OUTPUT NODEFVAL "eq53"
-- Retrieval info: USED_PORT: eq54 0 0 0 0 OUTPUT NODEFVAL "eq54"
-- Retrieval info: USED_PORT: eq55 0 0 0 0 OUTPUT NODEFVAL "eq55"
-- Retrieval info: USED_PORT: eq56 0 0 0 0 OUTPUT NODEFVAL "eq56"
-- Retrieval info: USED_PORT: eq57 0 0 0 0 OUTPUT NODEFVAL "eq57"
-- Retrieval info: USED_PORT: eq58 0 0 0 0 OUTPUT NODEFVAL "eq58"
-- Retrieval info: USED_PORT: eq59 0 0 0 0 OUTPUT NODEFVAL "eq59"
-- Retrieval info: USED_PORT: eq6 0 0 0 0 OUTPUT NODEFVAL "eq6"
-- Retrieval info: USED_PORT: eq60 0 0 0 0 OUTPUT NODEFVAL "eq60"
-- Retrieval info: USED_PORT: eq61 0 0 0 0 OUTPUT NODEFVAL "eq61"
-- Retrieval info: USED_PORT: eq62 0 0 0 0 OUTPUT NODEFVAL "eq62"
-- Retrieval info: USED_PORT: eq63 0 0 0 0 OUTPUT NODEFVAL "eq63"
-- Retrieval info: USED_PORT: eq64 0 0 0 0 OUTPUT NODEFVAL "eq64"
-- Retrieval info: USED_PORT: eq65 0 0 0 0 OUTPUT NODEFVAL "eq65"
-- Retrieval info: USED_PORT: eq66 0 0 0 0 OUTPUT NODEFVAL "eq66"
-- Retrieval info: USED_PORT: eq67 0 0 0 0 OUTPUT NODEFVAL "eq67"
-- Retrieval info: USED_PORT: eq68 0 0 0 0 OUTPUT NODEFVAL "eq68"
-- Retrieval info: USED_PORT: eq69 0 0 0 0 OUTPUT NODEFVAL "eq69"
-- Retrieval info: USED_PORT: eq7 0 0 0 0 OUTPUT NODEFVAL "eq7"
-- Retrieval info: USED_PORT: eq70 0 0 0 0 OUTPUT NODEFVAL "eq70"
-- Retrieval info: USED_PORT: eq8 0 0 0 0 OUTPUT NODEFVAL "eq8"
-- Retrieval info: USED_PORT: eq9 0 0 0 0 OUTPUT NODEFVAL "eq9"
-- Retrieval info: CONNECT: @data 0 0 8 0 data 0 0 8 0
-- Retrieval info: CONNECT: eq0 0 0 0 0 @eq 0 0 1 0
-- Retrieval info: CONNECT: eq1 0 0 0 0 @eq 0 0 1 1
-- Retrieval info: CONNECT: eq10 0 0 0 0 @eq 0 0 1 10
-- Retrieval info: CONNECT: eq11 0 0 0 0 @eq 0 0 1 11
-- Retrieval info: CONNECT: eq12 0 0 0 0 @eq 0 0 1 12
-- Retrieval info: CONNECT: eq13 0 0 0 0 @eq 0 0 1 13
-- Retrieval info: CONNECT: eq14 0 0 0 0 @eq 0 0 1 14
-- Retrieval info: CONNECT: eq15 0 0 0 0 @eq 0 0 1 15
-- Retrieval info: CONNECT: eq16 0 0 0 0 @eq 0 0 1 16
-- Retrieval info: CONNECT: eq17 0 0 0 0 @eq 0 0 1 17
-- Retrieval info: CONNECT: eq18 0 0 0 0 @eq 0 0 1 18
-- Retrieval info: CONNECT: eq19 0 0 0 0 @eq 0 0 1 19
-- Retrieval info: CONNECT: eq2 0 0 0 0 @eq 0 0 1 2
-- Retrieval info: CONNECT: eq20 0 0 0 0 @eq 0 0 1 20
-- Retrieval info: CONNECT: eq21 0 0 0 0 @eq 0 0 1 21
-- Retrieval info: CONNECT: eq22 0 0 0 0 @eq 0 0 1 22
-- Retrieval info: CONNECT: eq23 0 0 0 0 @eq 0 0 1 23
-- Retrieval info: CONNECT: eq24 0 0 0 0 @eq 0 0 1 24
-- Retrieval info: CONNECT: eq25 0 0 0 0 @eq 0 0 1 25
-- Retrieval info: CONNECT: eq26 0 0 0 0 @eq 0 0 1 26
-- Retrieval info: CONNECT: eq27 0 0 0 0 @eq 0 0 1 27
-- Retrieval info: CONNECT: eq28 0 0 0 0 @eq 0 0 1 28
-- Retrieval info: CONNECT: eq29 0 0 0 0 @eq 0 0 1 29
-- Retrieval info: CONNECT: eq3 0 0 0 0 @eq 0 0 1 3
-- Retrieval info: CONNECT: eq30 0 0 0 0 @eq 0 0 1 30
-- Retrieval info: CONNECT: eq31 0 0 0 0 @eq 0 0 1 31
-- Retrieval info: CONNECT: eq32 0 0 0 0 @eq 0 0 1 32
-- Retrieval info: CONNECT: eq33 0 0 0 0 @eq 0 0 1 33
-- Retrieval info: CONNECT: eq34 0 0 0 0 @eq 0 0 1 34
-- Retrieval info: CONNECT: eq35 0 0 0 0 @eq 0 0 1 35
-- Retrieval info: CONNECT: eq36 0 0 0 0 @eq 0 0 1 36
-- Retrieval info: CONNECT: eq37 0 0 0 0 @eq 0 0 1 37
-- Retrieval info: CONNECT: eq38 0 0 0 0 @eq 0 0 1 38
-- Retrieval info: CONNECT: eq39 0 0 0 0 @eq 0 0 1 39
-- Retrieval info: CONNECT: eq4 0 0 0 0 @eq 0 0 1 4
-- Retrieval info: CONNECT: eq40 0 0 0 0 @eq 0 0 1 40
-- Retrieval info: CONNECT: eq41 0 0 0 0 @eq 0 0 1 41
-- Retrieval info: CONNECT: eq42 0 0 0 0 @eq 0 0 1 42
-- Retrieval info: CONNECT: eq43 0 0 0 0 @eq 0 0 1 43
-- Retrieval info: CONNECT: eq44 0 0 0 0 @eq 0 0 1 44
-- Retrieval info: CONNECT: eq45 0 0 0 0 @eq 0 0 1 45
-- Retrieval info: CONNECT: eq46 0 0 0 0 @eq 0 0 1 46
-- Retrieval info: CONNECT: eq47 0 0 0 0 @eq 0 0 1 47
-- Retrieval info: CONNECT: eq48 0 0 0 0 @eq 0 0 1 48
-- Retrieval info: CONNECT: eq49 0 0 0 0 @eq 0 0 1 49
-- Retrieval info: CONNECT: eq5 0 0 0 0 @eq 0 0 1 5
-- Retrieval info: CONNECT: eq50 0 0 0 0 @eq 0 0 1 50
-- Retrieval info: CONNECT: eq51 0 0 0 0 @eq 0 0 1 51
-- Retrieval info: CONNECT: eq52 0 0 0 0 @eq 0 0 1 52
-- Retrieval info: CONNECT: eq53 0 0 0 0 @eq 0 0 1 53
-- Retrieval info: CONNECT: eq54 0 0 0 0 @eq 0 0 1 54
-- Retrieval info: CONNECT: eq55 0 0 0 0 @eq 0 0 1 55
-- Retrieval info: CONNECT: eq56 0 0 0 0 @eq 0 0 1 56
-- Retrieval info: CONNECT: eq57 0 0 0 0 @eq 0 0 1 57
-- Retrieval info: CONNECT: eq58 0 0 0 0 @eq 0 0 1 58
-- Retrieval info: CONNECT: eq59 0 0 0 0 @eq 0 0 1 59
-- Retrieval info: CONNECT: eq6 0 0 0 0 @eq 0 0 1 6
-- Retrieval info: CONNECT: eq60 0 0 0 0 @eq 0 0 1 60
-- Retrieval info: CONNECT: eq61 0 0 0 0 @eq 0 0 1 61
-- Retrieval info: CONNECT: eq62 0 0 0 0 @eq 0 0 1 62
-- Retrieval info: CONNECT: eq63 0 0 0 0 @eq 0 0 1 63
-- Retrieval info: CONNECT: eq64 0 0 0 0 @eq 0 0 1 64
-- Retrieval info: CONNECT: eq65 0 0 0 0 @eq 0 0 1 65
-- Retrieval info: CONNECT: eq66 0 0 0 0 @eq 0 0 1 66
-- Retrieval info: CONNECT: eq67 0 0 0 0 @eq 0 0 1 67
-- Retrieval info: CONNECT: eq68 0 0 0 0 @eq 0 0 1 68
-- Retrieval info: CONNECT: eq69 0 0 0 0 @eq 0 0 1 69
-- Retrieval info: CONNECT: eq7 0 0 0 0 @eq 0 0 1 7
-- Retrieval info: CONNECT: eq70 0 0 0 0 @eq 0 0 1 70
-- Retrieval info: CONNECT: eq8 0 0 0 0 @eq 0 0 1 8
-- Retrieval info: CONNECT: eq9 0 0 0 0 @eq 0 0 1 9
-- Retrieval info: GEN_FILE: TYPE_NORMAL decode.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL decode.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL decode.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL decode.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL decode_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
