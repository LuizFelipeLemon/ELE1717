    Mac OS X            	   2   �      �                                      ATTR       �   �   F                  �   F  com.apple.quarantine q/0001;56f1d3a7;Google\x20Chrome;0D0B0B7A-70C2-407F-A0D8-C567BDD98245 